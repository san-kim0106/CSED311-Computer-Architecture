module Memory #(parameter MEM_DEPTH = 16384) (input reset,
                                              input clk,
                                              input [31:0] addr,    // address of the memory
                                              input [31:0] din,     // data to be written
                                              input mem_read,       // control signal
                                              input mem_write,      // control signal
                                              output reg [31:0] dout);  // output of the data memory at addr
  integer i;
  // Memory
  reg [31:0] mem[0: MEM_DEPTH - 1];
  // Do not touch mem_addr
  wire [31:0] mem_addr;
  assign mem_addr = {2'b00, addr >> 2};

  // Asynchrnously read data from the memory
  always @(addr, mem_read) begin
    if (mem_read) begin
      dout = mem[mem_addr];
    end else begin
      dout = 32'b0;
    end
    // $display("addr: %d | mem_read: %d | dout: %d", addr, mem_read, dout); //! DEBUGGING
  end

  always @(posedge clk) begin
    // Initialize data memory (do not touch)
    if (reset) begin
      for (i = 0; i < MEM_DEPTH; i = i + 1)
        mem[i] = 32'b0;
      // Provide path of the file including instructions with binary format
      $readmemh("C:\\Users\\sany0\\OneDrive\\Desktop\\CSED311-Computer-Architecture\\Labs\\Lab3\\lab3_tb\\test.txt", mem);
    end

    // Synchronously write data to the memory
    else begin
      if (mem_write) // Do not write to x0 register
        mem[mem_addr] <= din;
    end
  end
endmodule